'timescale 1ns/ 1ps

module AND(
    input SW1,
    input SW2,
    output LED
);
and u1 (SW1, SW2, LED);
endmodule